-- DIG_IN.VHD (a peripheral for SCOMP)
-- This device reads 16 digital inputs and provides
-- that data to SCOMP.

LIBRARY IEEE;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE LPM.LPM_COMPONENTS.ALL;

ENTITY DIG_IN IS
  PORT(
    IO_ADDR     : IN    STD_LOGIC_VECTOR(10 DOWNTO 0);
	 IO_READ     : IN    STD_LOGIC;
    EXT_WIRES   : IN    STD_LOGIC_VECTOR(15 DOWNTO 0);
    IO_DATA     : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END DIG_IN;

ARCHITECTURE a OF DIG_IN IS
  SIGNAL CHIP_SELECT : STD_LOGIC;

  BEGIN

	 CHIP_SELECT <=
      '1' WHEN (IO_ADDR = "00000000000") AND (IO_READ = '1')
		ELSE '0';

	IO_DATA <=
		EXT_WIRES WHEN CHIP_SELECT = '1'
		ELSE "ZZZZZZZZZZZZZZZZ";
		
END a;

