LIBRARY IEEE;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE LPM.LPM_COMPONENTS.ALL;

ENTITY Math_Peripheral IS
    PORT (
        CLOCK,
        RESETN   : IN    STD_LOGIC;
        IO_ADDR  : IN    STD_LOGIC_VECTOR(10 DOWNTO 0);
        IO_READ  : IN    STD_LOGIC;
        IO_WRITE : IN    STD_LOGIC;
        IO_DATA  : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END Math_Peripheral;
ARCHITECTURE a OF Math_Peripheral IS

    -- Internal registers
    SIGNAL x1, x2    : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL Result   : STD_LOGIC_VECTOR(7 DOWNTO 0);

    SIGNAL IO_EN : STD_LOGIC;
    SIGNAL IO_OUT : STD_LOGIC_VECTOR(15 DOWNTO 0);

	Begin --GoFromHere
    
    IO_EN <= IO_READ OR IO_WRITE;

    PROCESS (CLOCK, RESETN)
    BEGIN
        IF RESETN = '0' THEN
            x1 <= (OTHERS => '0');
            x2 <= (OTHERS => '0');
            Result <= (OTHERS => '0');
        ELSIF RISING_EDGE(CLOCK) THEN
         IF (IO_WRITE = '1') THEN
            CASE IO_ADDR IS
                WHEN "00100100000" =>  -- 0x90 MULT
                    x1 <= IO_DATA(7 DOWNTO 4);
                    x2 <= IO_DATA(3 DOWNTO 0);
                    Result <= ("0000" & x1) * ("0000" & x2);

                WHEN "00100100001" =>  -- 0x91 DIV
                    x1 <= IO_DATA(7 DOWNTO 4);
                    x2 <= IO_DATA(3 DOWNTO 0);
                    IF x2 /= "0000" THEN
                        Result <= RE("0000" & x1) / ("0000" & x2);
                    ELSE
                        Result <= (OTHERS => '0');
                    END IF;

                WHEN "00100100010" =>  -- 0x92 MOD
                    x1 <= IO_DATA(7 DOWNTO 4);
                    x2 <= IO_DATA(3 DOWNTO 0);
                    IF x2 /= "0000" THEN
                        Result <= ("0000" & x1) MOD ("0000" & x2);
                    ELSE
                        Result <= (OTHERS => '0');
                    END IF;

                WHEN OTHERS =>
                    NULL;
            END CASE;
        END IF;
    END IF;
END PROCESS;

    IO_DATA <= IO_OUT WHEN IO_READ = '1' ELSE (OTHERS => 'Z');
End a;